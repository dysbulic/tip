* W:\odin\hat\hat_controller.sch

* Schematics Version 8.0 - July 1997
* Wed Nov 06 12:06:08 2002



** Analysis setup **
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "hat_controller.net"
.INC "hat_controller.als"


.probe


.END
